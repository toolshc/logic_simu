��  CCircuit��  CSerializeHack           ��  CPart�� 
 CTextLabel  � �     C      �  � � �     B      �  I � T     A                    ���  COR�� 	 CTerminal  ����     	 	        �          �  ����                          �  ���               �            ����           ��    �� 	 CLogicOut�   ��      	        �            �$�           ��    ��  CAND�  ����      	        �          �  ����                          �  ����     	          �            ����           ��    ��  @�U�              @          �  @�U�     
                     �  l���               �            T�l�           ��    �� 	 CRailThru�  x�       d                   �  |�                            z�         ����    ��  � x� �      
 d                   �  � |� �                            � z� �    #    ����    ��  ` xa �       d                   �  ` |a �                            \ zd �    &    ����    ��  @ xA �       d       @          �  @ |A �              @            < zD �    )    ����    �� 	 CInverter�  @ HA ]                           �  @ tA �              @            4 \L t    -      ��    ��  � � 1                            � �     0      ��    ��  � � 1     
                       � �     2      ��    ��  @ A 1                            8 H     4      ��    ��  CLogicIn�� 	 CLatchKey  �       6   �  1                                9    ����     5�7�  � �       :   �  � � 1     
                       � �     <    ����     5�7�  H X       =   �  ` a 1                            \ d     ?    ����                   ���  CWire  ` �a y       A��� 
 CCrossOver  ^ �d �        ` 0a �       A�D�  � �� �      D�  ��        ` ���      A�  ����       A�D�  � �� �        � �� y      
 A�D�  ��        �y       A�  @ �A y       A�D�  ��      D�  ��        0�       A�  ���      A�  ����       A�D�  � �� �        � 0� �      
 A�D�  ��        � �A�     
 A�  @ �A �       A�D�  ^ �d �      D�  � �� �      D�  ��        @ �A�      A�  @ 0A I       A�  @ 0a 1      A�  � 0� 1     
 A�  � 01                    �                                I            S      Y   V     L   ! !   J # $ $   B & ' '   N ) * *   - ] - . . X 0 0 ` 2 2 _ 4 4 ^ 9 9 ` < < _ ? ? ^ C & C Z ? F F K F M B I  F J G T # L H O   X ) O \ O W 9 R L S  R T [ < V V Q J  . Y Y E Y U Y P N  4 - ] C 2 T 0 O             �$s�        @     +        @            @    "V  (      �                 
         $@      �? V               �? V         
         $@      �? V               �? V                 @      �? s 