��  CCircuit��  CSerializeHack           ��  CPart�� 
 CTextLabel  9D    C      �  � �     B      �  Q \     A          H   H     ��� 	 CLogicOut�� 	 CTerminal  ����               �            ����           ��    ��  COR�  p���               �          �  p���               �          �  ����               �            �|��           ��    ��  CAND�  ���               �          �  �	                          �   1               �            �           ��    ��  ����                          �  ����                          �  ����               �            ����           ��    ��  H-I               �          �  X-Y               �          �  DPYQ               �            ,DD\           ��    ��  �p�q                          �  ����                          �  �x�y               �            �l��     #      ��    ��  ���               �          �  ���              @          �  �1�               �            ��     '      ��    �� 	 CRailThru�  � � -       d                   �  � � 1                            � � .    ,    ����    *��  � � -       d                   �  � � 1     
                       | � .    /    ����    *��  @ A -       d       @          �  @ A 1              @            < D .    2    ����    *��  � � -       d       @          �  � � 1              @            � � .    5    ����    *��  xy-       d                   �  xy1                            t|.    8    ����    *��  ()-       d       @          �  ()1              @            $,.    ;    ����    ��  � �               �          �  ��               �          �  ��	               �            ���     >      ��    ��  �@A     	          �          �  �PQ                          �  $H9I               �            <$T     B      ��    ��  � �!                          �  �0�1              @          �  �(�)     	          �            ��4     F      ��    ��  X�m�               �          �  X�m�               �          �  ����               �            l���     J      ��    ��  ���               �          �  ���              @          �  $�9�               �            �$�     N      ��    ��  ����                          �  ����              @          �  ����               �            ����     R      ��    ��  ���               �          �  ���                          �  $�9�               �            �$�     V      ��    ��  ($)9                             0$    Z      ��    ��  CLogicIn�� 	 CLatchKey  8H'      \   �  P$Q9                            LT$    _    ����     �� 	 CInverter�  (8)M       	                   �  (d)y              @            L4d    b      ��    ��  ����              @          �  ����                          �  ����               �            �|��     e      ��    ��  � $� 9                            � � $    i      ��    [�]�  � � '      j   �  � $� 9                            � � $    l    ����     `��  � 8� M       	                   �  � d� y              @            � L� d    n      ��    `��  @ 8A M       	                   �  @ dA y              @            4 LL d    q      ��    ��  @ $A 9                            8 H $    t      ��    [�]�  P ` '      u   �  h $i 9                            d l $    w    ����         H   H     ���  CWire  ����      y�  p�q       y�  0 q      y�  pPq�       y�  XPqQ      y�  I       y�  ��I       y��� 
 CCrossOver  &|,�      ��  &�,�      ��  &�,�      ��  &�,�        (x)�       y�  xy       y���  vl|t      ��  v||�      ��  v�|�      ��  v�|�      ��  v�|�        xPy	       y�  x�	      y�  � ��        y���  � �� �        � �� �       y���  &�,�      ��  v�|�        � ���      y���  &�,�      ��  &�,�        (�)       y�  � ��        y�  � p� �       y���  � �� �      ��  � �� �      ��  &�,�      ��  v�|�        � ���      y���  � �� �      ��  � l� t        � 0�        y�  ����       y�  ����      y�  �	      y�  X�       y�  0��      y���  v||�      ��  v�|�        x8y�       y���  &,,4      ��  &,$      ��  &l,t      ��  &|,�        (�)�       y���  v�|�        (���      y���  � ,� 4      ��  � � $      ��  � �� �      ��  � �� �      ��  � l� t        � �� �       y���  &|,�      ��  v||�        � ���      y�  �  � q       y���  � l� t      ��  � l� t      ��  &l,t      ��  vl|t        � p�q      y�  �x��       y�  ����      y�  @ �A        y���  v�|�      ��  v�|�      ��  v�|�      ��  v|$      ��  v,|4        x�yQ       y���  v�|�        (���      y���  &,$      ��  � � $      ��  � � $      ��  v|$        �  �!      y���  &,,4      ��  � ,� 4      ��  v,|4        � 0�1      y���  � |� �        � 8� �       y���  � �� �      ��  � �� �      ��  &�,�      ��  v�|�        � ���      y���  � �� �      ��  &�,�      ��  v�|�        � ���      y���  � � $        � �� 1       y�  � �� !       y�  @ xA �       y�  8H�I      y�  ���       y�  ����      y�  xP�Q      y�  �(�)     	 y�  �(�A      	 y�  8�Y�      y�  8�9�       y�  8�Y�      y�  8�9�       y���  � |� �      ��  � �� �        � x� �       y���  ~ |� �        � 8� �       y�  ����      y�  ����       y�  x���      y�  ����       y�  ����      y���  &�,�      ��  v�|�        � ���      y���  ~ |� �      ��  � |� �      ��  � |� �      ��  &|,�      ��  v||�        @ ���      y�  (8Q9      y�  P8y9      y�  � 8� 9      y�  � 8� 9      y�  @ 8i 9      y�  h 8� 9          H   H     �    H   H         H   H      z   }   {    z  �   �    |  �   �    �      �   ! ! ~ # � # $ � $ % % � ' � ' ( � ( ) ) � � , - -   � / 0 0   � 2 3 3   � 5 6 6   � 8 9 9   � ; < <   > � > ? � ? @ @ � B � B C � C D D � F � F G � G H H � J � J K � K L L � N � N O � O P P � R � R S � S T T � V � V W � W X X � Z Z  _ _  b Z b c c � e � e f � f g g � i i l l n i n o o � q t q r r � t t w w    |  { ~  ! } �  ? � � � � � � � � � c � � 8 � � � � � � � � � � � � �  � , � � � � � � � � �  � � � � � ; � / � � � � � � � � � � �  � � � � � 5 �   � @    � ) � � � � � � � � � � � � � � � � � � � ( � � � � � � � � � � � � � � � � � $ � � � � � � � � � � � # % � � ' � 2 � � � � � � � � � � � � � � � O � � � � � � � � � F � � � � � � � G � � � � � � � � � � � � R � � � � � � � S � � � � � � r � D � � > L � � C H � � B � K � P � J X � � � � � o � � � � � N T � � W � V g � � � � � � f � � � � � � � � � � � e b _ � n l � q w �             �$s�        @     +        @            @    "V  (      �h                
         $@      �? V               �? V         
         $@      �? V               �? V                 @      �? s 